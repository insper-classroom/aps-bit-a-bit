-- Elementos de Sistemas
-- FlipFlopJK.vhd

library ieee;
use ieee.std_logic_1164.all;

entity FlipFlopJK is
	port(
		clock:  in std_logic;
		J:      in std_logic;
		K:      in std_logic;
		q:      out std_logic:= '0';
		notq:   out std_logic:= '1'
	);
end entity;

architecture arch of FlipFlopJK is
	signal q_int: std_logic := '0';
	signal entries: std_logic_vector(1 downto 0);

begin
	entries <= J & K;
	process(clock)
	begin
		if rising_edge(clock) then
			case entries is
				when "00" => 
					null;
				when "01" =>
					q_int <= '0';
				when "10" =>
					q_int <= '1';
				when others =>
					q_int <= not(q_int);
			end case;
		end if;
	end process;
	q <= q_int;
	notq <= not(q_int);
end architecture;