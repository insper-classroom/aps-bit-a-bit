-- Elementos de Sistemas
-- by Luciano Soares
-- Register64.vhd

Library ieee;
use ieee.std_logic_1164.all;

entity Register64 is
	port(
		clock:   in STD_LOGIC;
		input:   in STD_LOGIC_VECTOR(63 downto 0);
		load:    in STD_LOGIC;
		output: out STD_LOGIC_VECTOR(63 downto 0)
	);
end entity;

architecture arch of Register64 is

	component Register32 is
		port(
			clock:   in STD_LOGIC;
			input:   in STD_LOGIC_VECTOR(31 downto 0);
			load:    in STD_LOGIC;
			output: out STD_LOGIC_VECTOR(31 downto 0)
      );
	end component;

begin
	gen_bytes: for i in 0 to 1 generate
    constant hi : integer := i*32 + 31;
    constant lo : integer := i*32;
	begin
    	u_reg: Register32
    		port map(
        		clock  => clock,
        		input  => input(hi downto lo),
        		load   => load,
        		output => output(hi downto lo)
    		);
	end generate;
end architecture;