-- Elementos de Sistemas
-- by Luciano Soares
-- HalfAdder.vhd

-- Implementa Half Adder

Library ieee;
use ieee.std_logic_1164.all;

entity HalfAdder is
	port(
		a,b:         in STD_LOGIC;
		soma,vaium: out STD_LOGIC
	);
end entity;

architecture rtl of HalfAdder is
begin
    soma <= a xor b;
    vaium <= a and b;
end architecture;