--
-- Elementos de Sistemas - Aula 5 - Logica Combinacional
-- Rafael . Corsi @ insper . edu . br 
--
-- Arquivo exemplo para acionar os LEDs e ler os bottoes
-- da placa DE0-CV utilizada no curso de elementos de 
-- sistemas do 3s da eng. da computacao

----------------------------
-- Bibliotecas ieee       --
----------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.all;

----------------------------
-- Entrada e saidas do bloco
----------------------------
entity TopLevel is
	port(
		SW      : in  std_logic_vector(9 downto 0);
		KEY     : in  std_logic_vector(3 downto 0);
		LEDR    : out std_logic_vector(9 downto 0);
		HEX0     : out std_logic_vector(6 downto 0); -- 7seg0
        HEX1     : out std_logic_vector(6 downto 0); -- 7seg0
        HEX2     : out std_logic_vector(6 downto 0);
		HEX3     : out std_logic_vector(6 downto 0)
	);
end entity;

----------------------------
-- Implementacao do bloco -- 
----------------------------
architecture rtl of TopLevel is


component FlipFlopD is
	port(
		clock:  in std_logic;
		d:      in std_logic;
		clear:  in std_logic;
		preset: in std_logic;
		q:     out std_logic
	);
end component;

component Ram8 is 
	port(
		clock:   in  STD_LOGIC;
		input:   in  STD_LOGIC_VECTOR(15 downto 0);
		load:    in  STD_LOGIC;
		address: in  STD_LOGIC_VECTOR( 2 downto 0);
		output:  out STD_LOGIC_VECTOR(15 downto 0)
	);
end component;

component PC is
  port(
    clock     : in  STD_LOGIC;
    increment : in  STD_LOGIC;
    load      : in  STD_LOGIC;
    reset     : in  STD_LOGIC;
    input     : in  STD_LOGIC_VECTOR(15 downto 0);
    output    : out STD_LOGIC_VECTOR(15 downto 0) 
  );
end component;

component sevenseg is
	port (
		bcd : in  STD_LOGIC_VECTOR(3 downto 0);
		leds: out STD_LOGIC_VECTOR(6 downto 0)
		);
end component;

--------------
-- signals
--------------

signal clock, clear, set : std_logic;
signal HexBF35: std_logic_vector(15 downto 0);
signal ad: std_logic_vector(2 downto 0);
signal outRam: std_logic_vector(15 downto 0);
signal outPC: std_logic_vector(15 downto 0);
signal numero: std_logic_vector(15 downto 0);

---------------
-- implementacao
---------------
begin

Clock <= not KEY(0); -- os botoes quando nao apertado vale 1
                     -- e apertado 0, essa logica inverte iss
clear <= not KEY(1);
set	<= not KEY(2);
--ad <= SW(2 downto 0);
HexBF35 <= x"BF35";
numero <= x"BC75";

-- u0 : FlipFlopD port map (
-- 		clock    => Clock,
-- 		d        => SW(0),
-- 		clear    => clear,
-- 		preset   => set,
-- 		q        => LEDR(0)
-- 	);		

-- u1: Ram8
-- 	port map(
-- 		clock => Clock,
-- 		input => HexBF35,
-- 		load => set,
-- 		address => ad,
-- 		output => outRam
-- 	);

pc0: PC
	port map(
		clock     => Clock,
		increment => SW(0),
		load      => set,
		reset     => SW(1),
		input     => numero,
		output    => outPC
	);

s0: sevenseg
	port map(
		bcd => outPC(3 downto 0),
		leds => HEX0
	);
s1: sevenseg
	port map(
		bcd => outPC(7 downto 4),
		leds => HEX1
	);

s2: sevenseg
	port map(
		bcd => outPC(11 downto 8),
		leds => HEX2
	);
s3: sevenseg
	port map(
		bcd => outPC(15 downto 12),
		leds => HEX3
	);



end rtl;
