--
-- Elementos de Sistemas - Aula 5 - Logica Combinacional
-- Rafael . Corsi @ insper . edu . br
--
-- Arquivo exemplo para acionar os LEDs e ler os bottoes
-- da placa DE0-CV utilizada no curso de elementos de
-- sistemas do 3s da eng. da computacao

----------------------------
-- Bibliotecas ieee       --
----------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.all;

----------------------------
-- Entrada e saidas do bloco
----------------------------
entity TopLevel is
	port(
		CLOCK_50 : in  std_logic;
		SW       : in  std_logic_vector(9 downto 0);
		LEDR     : out std_logic_vector(9 downto 0);
		HEX0     : out std_logic_vector(6 downto 0);
		HEX1     : out std_logic_vector(6 downto 0);
		HEX2     : out std_logic_vector(6 downto 0)
	);
end entity;

----------------------------
-- Implementacao do bloco --
----------------------------
architecture rtl of TopLevel is

component conceitoa is
	port(
		CLOCK_50 : in  std_logic;
		SW       : in  std_logic_vector(9 downto 0);
        HEX0     : out std_logic_vector(6 downto 0); -- 7seg0
        HEX1     : out std_logic_vector(6 downto 0); -- 7seg0
        HEX2     : out std_logic_vector(6 downto 0); -- 7seg0
		LEDR     : out std_logic_vector(9 downto 0)
	);
end component;
--------------
-- signals
--------------
signal bcd : std_logic_vector(3 downto 0);

---------------
-- implementacao
---------------
begin
	--LEDR(0) <= SW(0);
	--LEDR(0) <= not SW(0);
	--LEDR(0) <= SW(0) or SW(1);
	--LEDR<= "1111111111" when SW="1001101010" else "0000000000";
	HEX1 <= "1111111";
	HEX2 <= "1111111";
	bcd <= SW(3) & SW(2) & SW(1) & SW(0);
	with bcd select
		HEX0 <= 	"1000000" when "0000", --0
					"1111001" when "0001", --1
					"0100100" when "0010", --2
					"0110000" when "0011", --3
					"0011001" when "0100", --4
					"0010010" when "0101", --5
					"0000010" when "0110", --6
					"1111000" when "0111", --7
					"0000000" when "1000", --8
					"0010000" when "1001", --9
					"0001000" when "1010", --A
					"0000011" when "1011", --B
					"1000110" when "1100", --C
					"0100001" when "1101", --D
					"0000110" when "1110", --E
					"0001110" when "1111", --F
					"1111111" when others;	
end rtl;
